

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity project_tb is
end project_tb;

architecture projecttb of project_tb is
constant c_CLOCK_PERIOD         : time := 15 ns;
signal   tb_done                : std_logic;
signal   mem_address            : std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst                 : std_logic := '0';
signal   tb_start               : std_logic := '0';
signal   tb_clk                 : std_logic := '0';
signal   mem_o_data,mem_i_data  : std_logic_vector (7 downto 0);
signal   enable_wire            : std_logic;
signal   mem_we                 : std_logic;

--signal o_N : std_logic_vector(7 downto 0);
--signal o_stato     : std_logic_vector(4 downto 0);
--signal o_indirizzo : std_logic_vector(15 downto 0);
--signal o_scritto : std_logic_vector(15 downto 0);
--signal o_numRighe : std_logic_vector(7 downto 0);
--signal o_numColonne : std_logic_vector(7 downto 0);
--signal o_pixel : std_logic_vector(7 downto 0);
--signal o_numPixel : std_logic_vector(7 downto 0);
--signal o_delta : std_logic_vector(8 downto 0);
--signal o_shift : std_logic_vector(7 downto 0);
--signal o_max : std_logic_vector(7 downto 0);
--signal o_min : std_logic_vector(7 downto 0);
--signal o_value : std_logic_vector(15 downto 0);

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);


signal RAM: ram_type := (0 => std_logic_vector(to_unsigned(  2  , 8)), 
                         1 => std_logic_vector(to_unsigned(  2  , 8)), 
                         2 => std_logic_vector(to_unsigned(  46  , 8)),  
                         3 => std_logic_vector(to_unsigned(  131  , 8)), 
                         4 => std_logic_vector(to_unsigned(  62  , 8)), 
                         5 => std_logic_vector(to_unsigned(  89  , 8)), 
                         others => (others =>'0'));         
			 -- Expected Output  6 -> 0                         
			 -- Expected Output  7 -> 255                         
			 -- Expected Output  8 -> 64                         
			 -- Expected Output  9 -> 172                         

component project_reti_logiche is
port (
      i_clk         : in  std_logic;
      i_rst         : in  std_logic;
      i_start       : in  std_logic;
      i_data        : in  std_logic_vector(7 downto 0);
      o_address     : out std_logic_vector(15 downto 0);
      o_done        : out std_logic;
      o_en          : out std_logic;
      o_we          : out std_logic;
      o_data        : out std_logic_vector(7 downto 0)

      --o_N : out std_logic_vector(7 downto 0);
      --o_stato     : out std_logic_vector(4 downto 0);
      --o_indirizzo : out std_logic_vector(15 downto 0);
      --o_scritto : out std_logic_vector(15 downto 0);
      --o_numRighe : out std_logic_vector(7 downto 0);
      --o_numColonne : out std_logic_vector(7 downto 0);
      --o_pixel : out std_logic_vector(7 downto 0);
      --o_numPixel : out std_logic_vector(7 downto 0);
      --o_delta : out std_logic_vector(8 downto 0);
      --o_shift : out std_logic_vector(7 downto 0);
      --o_max : out std_logic_vector(7 downto 0);
      --o_min : out std_logic_vector(7 downto 0);
      --o_value : out std_logic_vector(15 downto 0)
      );
end component project_reti_logiche;


begin
UUT: project_reti_logiche
port map (
          i_clk      	=> tb_clk,
          i_rst      	=> tb_rst,
          i_start       => tb_start,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address,
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
          o_we 		=> mem_we,
          o_data    	=> mem_i_data
          --o_numRighe  => o_numRighe,
          --o_numColonne => o_numColonne,
          --o_pixel => o_pixel,
          --o_numPixel => o_numPixel,
          --o_delta => o_delta,
          --o_shift => o_shift,
          --o_max => o_max,
          --o_min => o_min,
          --o_indirizzo => o_indirizzo,
          --o_scritto => o_scritto,
          --o_value => o_value,
          --o_stato => o_stato,
          --o_N => o_N
          );

p_CLK_GEN : process is
begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
end process p_CLK_GEN;


MEM : process(tb_clk)
begin
    if tb_clk'event and tb_clk = '1' then
        if enable_wire = '1' then
            if mem_we = '1' then
                RAM(conv_integer(mem_address))  <= mem_i_data;
                mem_o_data                      <= mem_i_data after 1 ns;
            else
                mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
            end if;
        end if;
    end if;
end process;


test : process is
begin 
    wait for 100 ns;
    wait for c_CLOCK_PERIOD;
    tb_rst <= '1';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_rst <= '0';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_start <= '1';
    wait for c_CLOCK_PERIOD;
    wait until tb_done = '1';
    wait for c_CLOCK_PERIOD;
    tb_start <= '0';
    wait until tb_done = '0';
    wait for 100 ns;

    -- Immagine originale =  [46, 131, 62, 89]  
    -- Immagine di output =  [0, 255, 64, 172]  
    
    assert RAM(6) = std_logic_vector(to_unsigned( 0 , 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(6))))  severity failure;
    assert RAM(7) = std_logic_vector(to_unsigned( 255 , 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(7))))  severity failure;
    assert RAM(8) = std_logic_vector(to_unsigned( 64 , 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(8))))  severity failure;
    assert RAM(9) = std_logic_vector(to_unsigned( 172 , 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

    assert false report "Simulation Ended! TEST PASSATO" severity failure;
end process test;

end projecttb; 


